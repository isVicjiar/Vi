// Fetch file

module fetch(
input		clock,
input		reset,

output	[31:0]	instruction);

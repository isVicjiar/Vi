// Branch predictor

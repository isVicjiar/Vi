# Main module of the project

module vi_core (
# Core inputs
# Core outputs);

wire A;

register register(
	.clock		(),
	.reset		(),
	.write_enable	(),
	.write_addr	(),
);

// File for the bypass controller

module bypass_ctrl (
input clk_i,
input rsn_i,
input read_addr_a_i,
input read_addr_b_i,
input exe_data_i,
input exe_addr_i,
input exe_wr_en_i,
input mult1_data_i,
input mult1_addr_i,
input mult1_wr_en_i,
input mult2_data_i,
input mult2_addr_i,
input mult2_wr_en_i,
input mult3_data_i,
input mult3_addr_i,
input mult3_wr_en_i,
input mult4_data_i,
input mult4_addr_i,
input mult4_wr_en_i,
input mult5_data_i,
input mult5_addr_i,
input mult5_wr_en_i,
input cache_data_i,
input cache_addr_i,
input cache_wr_en_i,
input write_data_i,
input write_addr_i,
input write_en_i,
output bypass_a_en_o,
output bypass_b_en_o,
output bypass_data_a_o,
output bypass_data_b_o,
output stall_core_o
);
